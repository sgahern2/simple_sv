module sv_loops;
  initial begin
    repeat ();
  end


endmodule

